netcdf chirp_init {
dimensions:
        nfov = 9;
        nchan = 1679;
        nobs = 12150;
	utc_tuple = 8 ;
variables:
	float rad(nobs, nchan) ;
		string rad:units = "mW/(m2 sr cm-1)" ;
		string rad:ancillary_variables = "rad_lw_qc" ;
		string rad:long_name = "real spectral radiance" ;
		string rad:standard_name = "toa_outgoing_radiance_per_unit_wavenumber" ;
		string rad:coordinates = "lon lat" ;
		string rad:description = "real spectral radiance" ;
		rad:_FillValue = 9.96921e+36f ;
		string rad:coverage_content_type = "physicalMeasurement" ;

        byte rad_qc(nobs) ;
                string rad_qc:units = "1" ;
                rad_qc:valid_range = 0b, 2b ;
                string rad_qc:long_name = "rad QC summary flag" ;
                string rad_qc:standard_name = "toa_outgoing_radiance_per_unit_wavenumber status_flag" ;
                string rad_qc:coordinates = "lon lat" ;
                string rad_qc:description = "rad QC summary flag" ;
                rad_qc:_FillValue = -1b ;
                string rad_qc:coverage_content_type = "qualityInformation" ;
                string rad_qc:flag_meanings = "Best Good Do_Not_Use" ;
                rad_qc:flag_values = 0b, 1b, 2b ;

        byte chan_qc(nchan) ;
                string chan_qc:units = "1" ;
                chan_qc:valid_range = 0b, 2b ;
                string chan_qc:long_name = "rad synthetic fraction flag" ;
                string chan_qc:standard_name = "radiance synthetic fraction flag" ;
                string chan_qc:coordinates = "lon lat" ;
                string chan_qc:description = "rad synthetic fraction flag" ;
                chan_qc:_FillValue = -1b ;
                string chan_qc:coverage_content_type = "qualityInformation" ;
                string chan_qc:flag_meanings = "Best Good Do_Not_Use" ;
                chan_qc:flag_values = 0b, 1b, 2b ;

	float synfrac(nchan) ;
		string synfrac:units = "synthetic fraction (ratio)" ;
		string synfrac:long_name = "synthetic channel fraction" ;
		string synfrac:description = "synthetic channel fraction" ;
		synfrac:_FillValue = 9.96921e+36f ;
		string synfrac:coverage_content_type = "qualityInformation" ;

	float nedn(nfov, nchan) ;
		string nedn:units = "mW/(m2 sr cm-1)" ;
		string nedn:long_name = "noise equivalent differential radiance" ;
		string nedn:description = "noise equivalent differential radiance" ;
		nedn:_FillValue = 9.96921e+36f ;
		string nedn:coverage_content_type = "qualityInformation" ;

	double obs_time_tai93(nobs) ;
		string obs_time_tai93:units = "seconds since 1993-01-01 00:00" ;
		obs_time_tai93:valid_range = -2934835217., 3376598410. ;
		string obs_time_tai93:long_name = "earth view FOV midtime" ;
		string obs_time_tai93:standard_name = "time" ;
		string obs_time_tai93:description = "earth view observation midtime for each FOV" ;
		obs_time_tai93:_FillValue = 9.96920996838687e+36 ;
		string obs_time_tai93:coverage_content_type = "referenceInformation" ;
	ushort obs_time_utc(nobs, utc_tuple) ;
		string obs_time_utc:units = "1" ;
		string obs_time_utc:long_name = "earth view UTC FOV time" ;
		string obs_time_utc:coordinates = "utc_tuple_lbl" ;
		string obs_time_utc:description = "UTC earth view observation time as an array of integers: year, month, day, hour, minute, second, millisec, microsec" ;
		obs_time_utc:_FillValue = 65535US ;
		string obs_time_utc:coverage_content_type = "referenceInformation" ;
	float lat(nobs) ;
		string lat:units = "degrees_north" ;
		lat:valid_range = -90.f, 90.f ;
		string lat:long_name = "latitude" ;
		string lat:standard_name = "latitude" ;
		string lat:description = "latitude of FOV center" ;
		lat:_FillValue = 9.96921e+36f ;
		string lat:coverage_content_type = "referenceInformation" ;
		string lat:bounds = "lat_bnds" ;
	float lon(nobs) ;
		string lon:units = "degrees_east" ;
		lon:valid_range = -180.f, 180.f ;
		string lon:long_name = "longitude" ;
		string lon:standard_name = "longitude" ;
		string lon:description = "longitude of FOV center" ;
		lon:_FillValue = 9.96921e+36f ;
		string lon:coverage_content_type = "referenceInformation" ;
	float view_ang(nobs) ;
		string view_ang:units = "degree" ;
		view_ang:valid_range = 0.f, 180.f ;
		string view_ang:long_name = "view angle" ;
		string view_ang:standard_name = "sensor_view_angle" ;
		string view_ang:coordinates = "lon lat" ;
		string view_ang:description = "off nadir pointing angle" ;
		view_ang:_FillValue = 9.96921e+36f ;
		string view_ang:coverage_content_type = "referenceInformation" ;
	float sat_zen(nobs) ;
		string sat_zen:units = "degree" ;
		sat_zen:valid_range = 0.f, 180.f ;
		string sat_zen:long_name = "satellite zenith angle" ;
		string sat_zen:standard_name = "sensor_zenith_angle" ;
		string sat_zen:coordinates = "lon lat" ;
		string sat_zen:description = "satellite zenith angle at the center of the FOV" ;
		sat_zen:_FillValue = 9.96921e+36f ;
		string sat_zen:coverage_content_type = "referenceInformation" ;
	float sat_azi(nobs) ;
		string sat_azi:units = "degree" ;
		sat_azi:valid_range = 0.f, 360.f ;
		string sat_azi:long_name = "satellite azimuth angle" ;
		string sat_azi:standard_name = "sensor_azimuth_angle" ;
		string sat_azi:coordinates = "lon lat" ;
		string sat_azi:description = "satellite azimuth angle at the center of the FOV (clockwise from North)" ;
		sat_azi:_FillValue = 9.96921e+36f ;
		string sat_azi:coverage_content_type = "referenceInformation" ;
		string lon:bounds = "lon_bnds" ;
	float sol_zen(nobs) ;
		string sol_zen:units = "degree" ;
		sol_zen:valid_range = 0.f, 180.f ;
		string sol_zen:long_name = "solar zenith angle" ;
		string sol_zen:standard_name = "solar_zenith_angle" ;
		string sol_zen:coordinates = "lon lat" ;
		string sol_zen:description = "solar zenith angle at the center of the FOV" ;
		sol_zen:_FillValue = 9.96921e+36f ;
		string sol_zen:coverage_content_type = "referenceInformation" ;
	float sol_azi(nobs) ;
		string sol_azi:units = "degree" ;
		sol_azi:valid_range = 0.f, 360.f ;
		string sol_azi:long_name = "solar azimuth angle" ;
		string sol_azi:standard_name = "solar_azimuth_angle" ;
		string sol_azi:coordinates = "lon lat" ;
		string sol_azi:description = "solar azimuth angle at the center of the FOV (clockwise from North)" ;
		sol_azi:_FillValue = 9.96921e+36f ;
		string sol_azi:coverage_content_type = "referenceInformation" ;
	float land_frac(nobs) ;
		string land_frac:units = "1" ;
		land_frac:valid_range = 0.f, 1.f ;
		string land_frac:long_name = "land fraction" ;
		string land_frac:standard_name = "land_area_fraction" ;
		string land_frac:coordinates = "lon lat" ;
		string land_frac:description = "land fraction over the FOV" ;
		land_frac:_FillValue = 9.96921e+36f ;
		string land_frac:coverage_content_type = "referenceInformation" ;
		string land_frac:cell_methods = "area: mean (beam-weighted)" ;
	float surf_alt(nobs) ;
		string surf_alt:units = "m" ;
		string surf_alt:ancillary_variables = "surf_alt_sdev" ;
		surf_alt:valid_range = -500.f, 10000.f ;
		string surf_alt:long_name = "surface altitude" ;
		string surf_alt:standard_name = "surface_altitude" ;
		string surf_alt:coordinates = "lon lat" ;
		string surf_alt:description = "mean surface altitude wrt  earth model over the FOV" ;
		surf_alt:_FillValue = 9.96921e+36f ;
		string surf_alt:coverage_content_type = "referenceInformation" ;
		string surf_alt:cell_methods = "area: mean (beam-weighted)" ;
	float surf_alt_sdev(nobs) ;
		string surf_alt_sdev:units = "m" ;
		surf_alt_sdev:valid_range = 0.f, 10000.f ;
		string surf_alt_sdev:long_name = "surface altitude standard deviation" ;
		string surf_alt_sdev:coordinates = "lon lat" ;
		string surf_alt_sdev:description = "standard deviation of surface altitude within the FOV" ;
		surf_alt_sdev:_FillValue = 9.96921e+36f ;
		string surf_alt_sdev:coverage_content_type = "qualityInformation" ;
		string surf_alt_sdev:cell_methods = "area: standard_deviation (beam-weighted)" ;
	ubyte instrument_state(nobs) ;
		string instrument_state:units = "1" ;
		string instrument_state:long_name = "instrument state" ;
		string instrument_state:coordinates = "lon lat" ;
		string instrument_state:description = "instrument/data state: 0/\'Process\' - Data is usable for science; 1/\'Special\' - Observations are valid but instrument is not configured for science data (ex: stare mode); 2/\'Erroneous\' - Data is not usable (ex: checksum error); 3/\'Missing\' - No data was received." ;
		instrument_state:_FillValue = 255UB ;
		string instrument_state:coverage_content_type = "qualityInformation" ;
		string instrument_state:flag_meanings = "Process Special Erroneous Missing" ;
		instrument_state:flag_values = 0UB, 1UB, 2UB, 3UB ;

	float subsat_lat(nobs) ;
		string subsat_lat:units = "degrees_north" ;
		subsat_lat:valid_range = -90.f, 90.f ;
		string subsat_lat:long_name = "sub-satellite latitude" ;
		string subsat_lat:standard_name = "latitude" ;
		string subsat_lat:description = "sub-satellite latitude at scan_mid_time" ;
		subsat_lat:_FillValue = 9.96921e+36f ;
		string subsat_lat:coverage_content_type = "referenceInformation" ;
	float subsat_lon(nobs) ;
		string subsat_lon:units = "degrees_east" ;
		subsat_lon:valid_range = -180.f, 180.f ;
		string subsat_lon:long_name = "sub-satellite longitude" ;
		string subsat_lon:standard_name = "longitude" ;
		string subsat_lon:description = "sub-satellite longitude at scan_mid_time" ;
		subsat_lon:_FillValue = 9.96921e+36f ;
		string subsat_lon:coverage_content_type = "referenceInformation" ;
	double scan_mid_time(nobs) ;
		string scan_mid_time:units = "seconds since 1993-01-01 00:00" ;
		scan_mid_time:valid_range = -2934835217., 3376598410. ;
		string scan_mid_time:long_name = "midscan TAI93" ;
		string scan_mid_time:standard_name = "time" ;
		string scan_mid_time:coordinates = "subsat_lon subsat_lat" ;
		string scan_mid_time:description = "TAI93 at  middle of earth scene scans" ;
		scan_mid_time:_FillValue = 9.96920996838687e+36 ;
		string scan_mid_time:coverage_content_type = "referenceInformation" ;
	float sat_alt(nobs) ;
		string sat_alt:units = "m" ;
		sat_alt:valid_range = 100000.f, 1000000.f ;
		string sat_alt:long_name = "satellite altitude" ;
		string sat_alt:standard_name = "altitude" ;
		string sat_alt:coordinates = "subsat_lon subsat_lat" ;
		string sat_alt:description = "satellite altitude with respect to earth model at scan_mid_time" ;
		sat_alt:_FillValue = 9.96921e+36f ;
		string sat_alt:coverage_content_type = "referenceInformation" ;
	float sun_glint_lat(nobs) ;
		string sun_glint_lat:units = "degrees_north" ;
		sun_glint_lat:valid_range = -90.f, 90.f ;
		string sun_glint_lat:long_name = "sun glint latitude" ;
		string sun_glint_lat:standard_name = "latitude" ;
		string sun_glint_lat:coordinates = "subsat_lon subsat_lat" ;
		string sun_glint_lat:description = "sun glint spot latitude at scan_mid_time.  Fill for night observations." ;
		sun_glint_lat:_FillValue = 9.96921e+36f ;
		string sun_glint_lat:coverage_content_type = "referenceInformation" ;
	float sun_glint_lon(nobs) ;
		string sun_glint_lon:units = "degrees_east" ;
		sun_glint_lon:valid_range = -180.f, 180.f ;
		string sun_glint_lon:long_name = "sun glint longitude" ;
		string sun_glint_lon:standard_name = "longitude" ;
		string sun_glint_lon:coordinates = "subsat_lon subsat_lat" ;
		string sun_glint_lon:description = "sun glint spot longitude at scan_mid_time.  Fill for night observations." ;
		sun_glint_lon:_FillValue = 9.96921e+36f ;
		string sun_glint_lon:coverage_content_type = "referenceInformation" ;
	ubyte asc_flag(nobs) ;
		string asc_flag:units = "1" ;
		asc_flag:valid_range = 0UB, 1UB ;
		string asc_flag:long_name = "ascending orbit flag" ;
		string asc_flag:coordinates = "subsat_lon subsat_lat" ;
		string asc_flag:description = "ascending orbit flag: 1 if ascending, 0 descending" ;
		asc_flag:_FillValue = 255UB ;
		string asc_flag:coverage_content_type = "referenceInformation" ;
		string asc_flag:flag_meanings = "descending ascending" ;
		asc_flag:flag_values = 0UB, 1UB ;

	ubyte airs_xtrack(nobs) ;
		string airs_xtrack:units = "1" ;
		airs_xtrack:valid_range = 1UB, 90UB ;
		string airs_xtrack:long_name = "field of regard number" ;
		string airs_xtrack:description = "field of regard number" ;
		airs_xtrack:_FillValue = 255UB ;
		string airs_xtrack:coverage_content_type = "auxiliaryInformation" ;

	ubyte airs_atrack(nobs) ;
		string airs_atrack:units = "1" ;
		airs_atrack:valid_range = 1UB, 135UB ;
		string airs_atrack:long_name = "field of view number" ;
		string airs_atrack:description = "field of view number" ;
		airs_atrack:_FillValue = 255UB ;
		string airs_atrack:coverage_content_type = "auxiliaryInformation" ;

	ubyte fov(nobs) ;
		string fov:units = "1" ;
		fov:valid_range = 1UB, 9UB ;
		string fov:long_name = "field of view number" ;
		string fov:description = "field of view number" ;
		fov:_FillValue = 255UB ;
		string fov:coverage_content_type = "auxiliaryInformation" ;

	ubyte xtrack(nobs) ;
		string xtrack:units = "1" ;
		xtrack:valid_range = 1UB, 30UB ;
		string xtrack:long_name = "field of regard number" ;
		string xtrack:description = "field of regard number" ;
		xtrack:_FillValue = 255UB ;
		string xtrack:coverage_content_type = "auxiliaryInformation" ;

	ubyte atrack(nobs) ;
		string xtrack:units = "1" ;
		xtrack:valid_range = 1UB, 45UB ;
		string xtrack:long_name = "scan index" ;
		string xtrack:description = "scan index" ;
		xtrack:_FillValue = 255UB ;
		string xtrack:coverage_content_type = "auxiliaryInformation" ;

	double wnum(nchan) ;
		string wnum:units = "cm-1" ;
		wnum:valid_range = 648.75, 2555.0 ;
		string wnum:long_name = "longwave wavenumber" ;
		string wnum:standard_name = "sensor_band_central_radiation_wavenumber" ;
		string wnum:description = "longwave wavenumber" ;
		wnum:_FillValue = 9.96920996838687e+36 ;
		string wnum:coverage_content_type = "auxiliaryInformation" ;

// global attributes:
		string :keywords = "EARTH SCIENCE > SPECTRAL/ENGINEERING > INFRARED WAVELENGTHS > INFRARED RADIANCE" ;
		string :processing_level = "1C" ;
		string :comment = "" ;
		string :acknowledgment = "Support for this research was provided by NASA." ;
		string :references = "" ;
		string :contributor_name = "UMBC Atmospheric Spectroscopy Laboratory: Larrabee Strow" ;
		string :contributor_role = "CrIS L1B Scientist" ;
		:license = "Freely Distributed" ;
		:product_name = "CHIRP" ;
		:product_name_version = "01a" ;
}

