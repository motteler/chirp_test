netcdf chirp_1330 {
dimensions:
	fov = 9 ;
	obs = 12150 ;
	wnum = 1679 ;
	fov_poly = 8 ;
	utc_tuple = 8 ;
variables:
	string obs_id(obs) ;
		string obs_id:long_name = "observation id" ;
		string obs_id:coverage_content_type = "referenceInformation" ;
		string obs_id:description = "unique earth view observation identifier." ;
	double obs_time_tai93(obs) ;
		obs_time_tai93:valid_range = -2934835217., 3376598410. ;
		string obs_time_tai93:long_name = "earth view FOV midtime" ;
		obs_time_tai93:_FillValue = 9.96920996838687e+36 ;
		string obs_time_tai93:coverage_content_type = "referenceInformation" ;
		string obs_time_tai93:standard_name = "time" ;
		string obs_time_tai93:units = "seconds since 1993-01-01 00:00" ;
		string obs_time_tai93:description = "earth view observation midtime for each FOV" ;
		string obs_time_tai93:AIRS_HDF_name = "Time" ;
	ushort obs_time_utc(obs, utc_tuple) ;
		string obs_time_utc:long_name = "earth view UTC FOV time" ;
		string obs_time_utc:coordinates = "utc_tuple_lbl" ;
		obs_time_utc:_FillValue = 65535US ;
		string obs_time_utc:coverage_content_type = "referenceInformation" ;
		string obs_time_utc:description = "UTC earth view observation time as an array of integers: year, month, day, hour, minute, second, millisec, microsec" ;
	float lat(obs) ;
		lat:valid_range = -90.f, 90.f ;
		string lat:long_name = "latitude" ;
		lat:_FillValue = 9.96921e+36f ;
		string lat:bounds = "lat_bnds" ;
		string lat:coverage_content_type = "referenceInformation" ;
		string lat:standard_name = "latitude" ;
		string lat:units = "degrees_north" ;
		string lat:description = "latitude of FOV center" ;
		string lat:AIRS_HDF_name = "Latitude" ;
	float lon(obs) ;
		lon:valid_range = -180.f, 180.f ;
		string lon:long_name = "FOV longitude" ;
		lon:_FillValue = 9.96921e+36f ;
		string lon:bounds = "lon_bnds" ;
		string lon:coverage_content_type = "referenceInformation" ;
		string lon:standard_name = "longitude" ;
		string lon:units = "degrees_east" ;
		string lon:description = "longitude of FOV center" ;
		string lon:AIRS_HDF_name = "Longitude" ;
	float lat_bnds(obs, fov_poly) ;
		lat_bnds:valid_range = -90.f, 90.f ;
		string lat_bnds:long_name = "FOV boundary latitudes" ;
		lat_bnds:_FillValue = 9.96921e+36f ;
		string lat_bnds:coverage_content_type = "referenceInformation" ;
		string lat_bnds:units = "degrees_north" ;
		string lat_bnds:description = "latitudes of points forming a polygon around the perimeter of the FOV" ;
	float lon_bnds(obs, fov_poly) ;
		lon_bnds:valid_range = -180.f, 180.f ;
		string lon_bnds:long_name = "FOV boundary longitudes" ;
		lon_bnds:_FillValue = 9.96921e+36f ;
		string lon_bnds:coverage_content_type = "referenceInformation" ;
		string lon_bnds:units = "degrees_east" ;
		string lon_bnds:description = "longitudes of points forming a polygon around the perimeter of the FOV" ;
	float land_frac(obs) ;
		land_frac:valid_range = 0.f, 1.f ;
		string land_frac:long_name = "land fraction" ;
		string land_frac:coordinates = "lon lat" ;
		land_frac:_FillValue = 9.96921e+36f ;
		string land_frac:coverage_content_type = "referenceInformation" ;
		string land_frac:standard_name = "land_area_fraction" ;
		string land_frac:units = "1" ;
		string land_frac:description = "land fraction over the FOV" ;
		string land_frac:AIRS_HDF_name = "landFrac" ;
		string land_frac:cell_methods = "area: mean (beam-weighted)" ;
	float surf_alt(obs) ;
		string surf_alt:ancillary_variables = "surf_alt_sdev" ;
		surf_alt:valid_range = -500.f, 10000.f ;
		string surf_alt:long_name = "surface altitude" ;
		string surf_alt:coordinates = "lon lat" ;
		surf_alt:_FillValue = 9.96921e+36f ;
		string surf_alt:coverage_content_type = "referenceInformation" ;
		string surf_alt:standard_name = "surface_altitude" ;
		string surf_alt:units = "m" ;
		string surf_alt:description = "mean surface altitude wrt  earth model over the FOV" ;
		string surf_alt:AIRS_HDF_name = "topog" ;
		string surf_alt:cell_methods = "area: mean (beam-weighted)" ;
	float surf_alt_sdev(obs) ;
		surf_alt_sdev:valid_range = 0.f, 10000.f ;
		string surf_alt_sdev:long_name = "surface altitude standard deviation" ;
		string surf_alt_sdev:coordinates = "lon lat" ;
		surf_alt_sdev:_FillValue = 9.96921e+36f ;
		string surf_alt_sdev:coverage_content_type = "qualityInformation" ;
		string surf_alt_sdev:units = "m" ;
		string surf_alt_sdev:description = "standard deviation of surface altitude within the FOV" ;
		string surf_alt_sdev:AIRS_HDF_name = "topog_err" ;
		string surf_alt_sdev:cell_methods = "area: standard_deviation (beam-weighted)" ;
	float sun_glint_lat(obs) ;
		sun_glint_lat:valid_range = -90.f, 90.f ;
		string sun_glint_lat:long_name = "sun glint latitude" ;
		string sun_glint_lat:coordinates = "subsat_lon subsat_lat" ;
		sun_glint_lat:_FillValue = 9.96921e+36f ;
		string sun_glint_lat:coverage_content_type = "referenceInformation" ;
		string sun_glint_lat:standard_name = "latitude" ;
		string sun_glint_lat:units = "degrees_north" ;
		string sun_glint_lat:description = "sun glint spot latitude at scan_mid_time.  Fill for night observations." ;
		string sun_glint_lat:AIRS_HDF_name = "glintlat" ;
	float sun_glint_lon(obs) ;
		sun_glint_lon:valid_range = -180.f, 180.f ;
		string sun_glint_lon:long_name = "sun glint longitude" ;
		string sun_glint_lon:coordinates = "subsat_lon subsat_lat" ;
		sun_glint_lon:_FillValue = 9.96921e+36f ;
		string sun_glint_lon:coverage_content_type = "referenceInformation" ;
		string sun_glint_lon:standard_name = "longitude" ;
		string sun_glint_lon:units = "degrees_east" ;
		string sun_glint_lon:description = "sun glint spot longitude at scan_mid_time.  Fill for night observations." ;
		string sun_glint_lon:AIRS_HDF_name = "glintlon" ;
	float sol_zen(obs) ;
		sol_zen:valid_range = 0.f, 180.f ;
		string sol_zen:long_name = "solar zenith angle" ;
		string sol_zen:coordinates = "lon lat" ;
		sol_zen:_FillValue = 9.96921e+36f ;
		string sol_zen:coverage_content_type = "referenceInformation" ;
		string sol_zen:standard_name = "solar_zenith_angle" ;
		string sol_zen:units = "degree" ;
		string sol_zen:description = "solar zenith angle at the center of the FOV" ;
		string sol_zen:AIRS_HDF_name = "solzen" ;
	float sol_azi(obs) ;
		sol_azi:valid_range = 0.f, 360.f ;
		string sol_azi:long_name = "solar azimuth angle" ;
		string sol_azi:coordinates = "lon lat" ;
		sol_azi:_FillValue = 9.96921e+36f ;
		string sol_azi:coverage_content_type = "referenceInformation" ;
		string sol_azi:standard_name = "solar_azimuth_angle" ;
		string sol_azi:units = "degree" ;
		string sol_azi:description = "solar azimuth angle at the center of the FOV (clockwise from North)" ;
		string sol_azi:AIRS_HDF_name = "solazi" ;
	float sun_glint_dist(obs) ;
		sun_glint_dist:valid_range = 0.f, 3.e+07f ;
		string sun_glint_dist:long_name = "sun glint distance" ;
		string sun_glint_dist:coordinates = "lon lat" ;
		sun_glint_dist:_FillValue = 9.96921e+36f ;
		string sun_glint_dist:coverage_content_type = "referenceInformation" ;
		string sun_glint_dist:units = "m" ;
		string sun_glint_dist:description = "distance of sun glint spot to the center of the FOV" ;
		string sun_glint_dist:AIRS_HDF_name = "sun_glint_distance" ;
	float view_ang(obs) ;
		view_ang:valid_range = 0.f, 180.f ;
		string view_ang:long_name = "view angle" ;
		string view_ang:coordinates = "lon lat" ;
		view_ang:_FillValue = 9.96921e+36f ;
		string view_ang:coverage_content_type = "referenceInformation" ;
		string view_ang:standard_name = "sensor_view_angle" ;
		string view_ang:units = "degree" ;
		string view_ang:description = "off nadir pointing angle" ;
		string view_ang:AIRS_HDF_name = "scanang" ;
	float sat_zen(obs) ;
		sat_zen:valid_range = 0.f, 180.f ;
		string sat_zen:long_name = "satellite zenith angle" ;
		string sat_zen:coordinates = "lon lat" ;
		sat_zen:_FillValue = 9.96921e+36f ;
		string sat_zen:coverage_content_type = "referenceInformation" ;
		string sat_zen:standard_name = "sensor_zenith_angle" ;
		string sat_zen:units = "degree" ;
		string sat_zen:description = "satellite zenith angle at the center of the FOV" ;
		string sat_zen:AIRS_HDF_name = "satzen" ;
	float sat_azi(obs) ;
		sat_azi:valid_range = 0.f, 360.f ;
		string sat_azi:long_name = "satellite azimuth angle" ;
		string sat_azi:coordinates = "lon lat" ;
		sat_azi:_FillValue = 9.96921e+36f ;
		string sat_azi:coverage_content_type = "referenceInformation" ;
		string sat_azi:standard_name = "sensor_azimuth_angle" ;
		string sat_azi:units = "degree" ;
		string sat_azi:description = "satellite azimuth angle at the center of the FOV (clockwise from North)" ;
		string sat_azi:AIRS_HDF_name = "satazi" ;
	float sat_range(obs) ;
		sat_range:valid_range = 100000.f, 1.e+07f ;
		string sat_range:long_name = "satellite range" ;
		string sat_range:coordinates = "lon lat" ;
		sat_range:_FillValue = 9.96921e+36f ;
		string sat_range:coverage_content_type = "referenceInformation" ;
		string sat_range:units = "m" ;
		string sat_range:description = "line of sight distance between satellite and FOV center" ;
	ubyte asc_flag(obs) ;
		asc_flag:valid_range = 0UB, 1UB ;
		string asc_flag:long_name = "ascending orbit flag" ;
		string asc_flag:coordinates = "subsat_lon subsat_lat" ;
		asc_flag:_FillValue = 255UB ;
		asc_flag:flag_values = 0UB, 1UB ;
		string asc_flag:coverage_content_type = "referenceInformation" ;
		string asc_flag:description = "ascending orbit flag: 1 if ascending, 0 descending" ;
		string asc_flag:AIRS_HDF_name = "scan_node_type" ;
		string asc_flag:flag_meanings = "descending ascending" ;
	float subsat_lat(obs) ;
		subsat_lat:valid_range = -90.f, 90.f ;
		string subsat_lat:long_name = "sub-satellite latitude" ;
		subsat_lat:_FillValue = 9.96921e+36f ;
		string subsat_lat:coverage_content_type = "referenceInformation" ;
		string subsat_lat:standard_name = "latitude" ;
		string subsat_lat:units = "degrees_north" ;
		string subsat_lat:description = "sub-satellite latitude at scan_mid_time" ;
		string subsat_lat:AIRS_HDF_name = "sat_lat" ;
	float subsat_lon(obs) ;
		subsat_lon:valid_range = -180.f, 180.f ;
		string subsat_lon:long_name = "sub-satellite longitude" ;
		subsat_lon:_FillValue = 9.96921e+36f ;
		string subsat_lon:coverage_content_type = "referenceInformation" ;
		string subsat_lon:standard_name = "longitude" ;
		string subsat_lon:units = "degrees_east" ;
		string subsat_lon:description = "sub-satellite longitude at scan_mid_time" ;
		string subsat_lon:AIRS_HDF_name = "sat_lon" ;
	double scan_mid_time(obs) ;
		scan_mid_time:valid_range = -2934835217., 3376598410. ;
		string scan_mid_time:long_name = "midscan TAI93" ;
		string scan_mid_time:coordinates = "subsat_lon subsat_lat" ;
		scan_mid_time:_FillValue = 9.96920996838687e+36 ;
		string scan_mid_time:coverage_content_type = "referenceInformation" ;
		string scan_mid_time:standard_name = "time" ;
		string scan_mid_time:units = "seconds since 1993-01-01 00:00" ;
		string scan_mid_time:description = "TAI93 at  middle of earth scene scans" ;
		string scan_mid_time:AIRS_HDF_name = "nadirTAI" ;
	float sat_alt(obs) ;
		sat_alt:valid_range = 100000.f, 1000000.f ;
		string sat_alt:long_name = "satellite altitude" ;
		string sat_alt:coordinates = "subsat_lon subsat_lat" ;
		sat_alt:_FillValue = 9.96921e+36f ;
		string sat_alt:coverage_content_type = "referenceInformation" ;
		string sat_alt:standard_name = "altitude" ;
		string sat_alt:units = "m" ;
		string sat_alt:description = "satellite altitude with respect to earth model at scan_mid_time" ;
		string sat_alt:AIRS_HDF_name = "satheight" ;
	float local_solar_time(obs) ;
		local_solar_time:valid_range = 0.f, 24.f ;
		string local_solar_time:long_name = "local apparent solar time" ;
		string local_solar_time:coordinates = "lon lat" ;
		local_solar_time:_FillValue = 9.96921e+36f ;
		string local_solar_time:coverage_content_type = "referenceInformation" ;
		string local_solar_time:units = "hours" ;
		string local_solar_time:description = "local apparent solar time in hours from midnight" ;
	string utc_tuple_lbl(utc_tuple) ;
		string utc_tuple_lbl:long_name = "UTC date/time parts" ;
		string utc_tuple_lbl:coverage_content_type = "auxiliaryInformation" ;
		string utc_tuple_lbl:description = "names of the elements of UTC when it is expressed as an array of integers year,month,day,hour,minute,second,millisecond,microsecond" ;
	float rad(obs, wnum) ;
		string rad:units = "mW/(m2 sr cm-1)" ;
		string rad:ancillary_variables = "rad_qc synth_frac chan_qc" ;
		string rad:long_name = "spectral radiance" ;
		string rad:standard_name = "toa_outgoing_radiance_per_unit_wavenumber" ;
		string rad:coordinates = "lon lat" ;
		string rad:description = "spectral radiance" ;
		rad:_FillValue = 9.96921e+36f ;
		string rad:coverage_content_type = "physicalMeasurement" ;
	byte rad_qc(obs) ;
		rad_qc:valid_range = 0b, 2b ;
		string rad_qc:long_name = "rad QC" ;
		string rad_qc:standard_name = "toa_outgoing_radiance_per_unit_wavenumber status_flag" ;
		string rad_qc:coordinates = "lon lat" ;
		string rad_qc:description = "rad QC flag" ;
		rad_qc:_FillValue = -1b ;
		string rad_qc:coverage_content_type = "qualityInformation" ;
		string rad_qc:flag_meanings = "Best Good Do_Not_Use" ;
		rad_qc:flag_values = 0b, 1b, 2b ;
	float synth_frac(wnum) ;
		string synth_frac:units = "1" ;
		synth_frac:valid_range = 0.f, 1.f ;
		string synth_frac:long_name = "Fraction synthesized" ;
		string synth_frac:description = "File mean fraction of signal that is attributed to synthesized AIRS Level-1C values" ;
		synth_frac:_FillValue = 9.96921e+36f ;
		string synth_frac:coverage_content_type = "qualityInformation" ;
	byte chan_qc(wnum) ;
		chan_qc:valid_range = 0b, 2b ;
		string chan_qc:long_name = "Channel QC" ;
		string chan_qc:standard_name = "toa_outgoing_radiance_per_unit_wavenumber status_flag" ;
		string chan_qc:description = "Quality of each channel." ;
		chan_qc:_FillValue = -1b ;
		string chan_qc:coverage_content_type = "qualityInformation" ;
		string chan_qc:flag_meanings = "Best Good Do_Not_Use" ;
		chan_qc:flag_values = 0b, 1b, 2b ;
	float nedn(fov, wnum) ;
		string nedn:units = "mW/(m2 sr cm-1)" ;
		string nedn:long_name = "noise equivalent differential radiance" ;
		string nedn:description = "noise equivalent differential radiance" ;
		nedn:_FillValue = 9.96921e+36f ;
		string nedn:coverage_content_type = "qualityInformation" ;
	ubyte atrack(obs) ;
		string atrack:units = "1" ;
		atrack:valid_range = 1UB, 45UB ;
		string atrack:long_name = "Along-track FOR index" ;
		string atrack:coordinates = "lon lat" ;
		string atrack:axis = "Y" ;
		string atrack:description = "Along-track index of Field Of Regard" ;
		atrack:_FillValue = 255UB ;
		string atrack:coverage_content_type = "auxiliaryInformation" ;
	ubyte xtrack(obs) ;
		string xtrack:units = "1" ;
		xtrack:valid_range = 1UB, 30UB ;
		string xtrack:long_name = "Cross-track FOR index" ;
		string xtrack:coordinates = "lon lat" ;
		string xtrack:axis = "X" ;
		string xtrack:description = "Cross-track index of Field Of Regard" ;
		xtrack:_FillValue = 255UB ;
		string xtrack:coverage_content_type = "auxiliaryInformation" ;
	ubyte fov_num(obs) ;
		string fov_num:units = "1" ;
		fov_num:valid_range = 1UB, 9UB ;
		string fov_num:long_name = "Field Of View number" ;
		string fov_num:coordinates = "lon lat" ;
		string fov_num:description = "Field Of View number in FOR" ;
		fov_num:_FillValue = 255UB ;
		string fov_num:coverage_content_type = "auxiliaryInformation" ;
	ubyte airs_atrack(obs) ;
		string airs_atrack:units = "1" ;
		airs_atrack:valid_range = 1UB, 135UB ;
		string airs_atrack:long_name = "Along-track AIRS FOV index" ;
		string airs_atrack:coordinates = "lon lat" ;
		string airs_atrack:axis = "Y" ;
		string airs_atrack:description = "AIRS-like along-track index of Field Of View" ;
		airs_atrack:_FillValue = 255UB ;
		string airs_atrack:coverage_content_type = "auxiliaryInformation" ;
	ubyte airs_xtrack(obs) ;
		string airs_xtrack:units = "1" ;
		airs_xtrack:valid_range = 1UB, 90UB ;
		string airs_xtrack:long_name = "Cross-track AIRS FOV index" ;
		string airs_xtrack:coordinates = "lon lat" ;
		string airs_xtrack:axis = "X" ;
		string airs_xtrack:description = "AIRS-like cross-track index of Field Of View" ;
		airs_xtrack:_FillValue = 255UB ;
		string airs_xtrack:coverage_content_type = "auxiliaryInformation" ;
	double wnum(wnum) ;
		string wnum:units = "cm-1" ;
		wnum:valid_range = 640., 2700. ;
		string wnum:long_name = "wavenumber" ;
		string wnum:standard_name = "sensor_band_central_radiation_wavenumber" ;
		string wnum:description = "wavenumber" ;
		wnum:_FillValue = 9.96920996838687e+36 ;
		string wnum:coverage_content_type = "auxiliaryInformation" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.8.19" ;
		string :keywords = "EARTH SCIENCE > SPECTRAL/ENGINEERING > INFRARED WAVELENGTHS > INFRARED RADIANCE" ;
		string :Conventions = "CF-1.6, ACDD-1.3" ;
		string :history = "" ;
		string :source = "AIRS and CrIS instrument telemetry" ;
		string :processing_level = "1" ;
		string :product_name_type_id = "L1" ;
		string :comment = "" ;
		string :acknowledgment = "Support for this research was provided by NASA." ;
		string :license = "Limited to Sounder SIPS affiliates" ;
		string :standard_name_vocabulary = "CF Standard Name Table v28" ;
		string :date_created = "Unassigned" ;
		string :creator_name = "Unassigned" ;
		string :creator_email = "Unassigned" ;
		string :creator_url = "Unassigned" ;
		string :institution = "Unassigned" ;
		string :project = "Sounder SIPS" ;
		string :product_name_project = "SNDR" ;
		string :publisher_name = "Unassigned" ;
		string :publisher_email = "Unassigned" ;
		string :publisher_url = "Unassigned" ;
		string :geospatial_bounds = "" ;
		string :geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_lat_min = 9.96921e+36f ;
		:geospatial_lat_max = 9.96921e+36f ;
		:geospatial_lon_min = 9.96921e+36f ;
		:geospatial_lon_max = 9.96921e+36f ;
		string :time_coverage_start = "" ;
		string :time_of_first_valid_obs = "" ;
		string :time_coverage_mid = "" ;
		string :time_coverage_end = "" ;
		string :time_of_last_valid_obs = "" ;
		string :time_coverage_duration = "P0000-00-00T00:06:00" ;
		string :product_name_duration = "m06" ;
		string :creator_type = "institution" ;
		string :creator_institution = "Jet Propulsion Laboratory -- California Institute of Technology" ;
		string :product_version = "v01.00.00" ;
		string :keywords_vocabulary = "GCMD:GCMD Keywords" ;
		string :platform = "JPSS-1 > Joint Polar Satellite System - 1, SUOMI-NPP > Suomi National Polar-orbiting Partnership, AQUA > Earth Observing System" ;
		string :platform_vocabulary = "GCMD:GCMD Keywords" ;
		string :product_name_platform = "SSYN1330" ;
		string :instrument = "AIRS > Atmospheric Infrared Sounder, CrIS > Cross-track Infrared Sounder" ;
		string :instrument_vocabulary = "GCMD:GCMD Keywords" ;
		string :product_name_instr = "CHIRP" ;
		string :product_name = "" ;
		string :product_name_variant = "std" ;
		string :product_name_version = "vxx_xx_xx" ;
		string :product_name_producer = "T" ;
		string :product_name_timestamp = "yymmddhhmmss" ;
		string :product_name_extension = "nc" ;
		:granule_number = 0US ;
		string :product_name_granule_number = "g000" ;
		string :gran_id = "yyyymmddThhmm" ;
		:geospatial_lat_mid = 9.96921e+36f ;
		:geospatial_lon_mid = 9.96921e+36f ;
		string :featureType = "trajectory" ;
		string :data_structure = "trajectory" ;
		string :cdm_data_type = "Trajectory" ;
		string :id = "Unassigned" ;
		string :naming_authority = "Unassigned" ;
		string :identifier_product_doi = "Unassigned" ;
		string :identifier_product_doi_authority = "Unassigned" ;
		string :algorithm_version = "" ;
		string :production_host = "" ;
		string :format_version = "v02.01.15" ;
		string :input_file_names = "" ;
		string :input_file_types = "" ;
		string :input_file_dates = "" ;
		string :orbitDirection = "NA" ;
		string :day_night_flag = "NA" ;
		string :AutomaticQualityFlag = "Missing" ;
		string :AutomaticQualityFlagExplanation = "\'Passed\': all spectra are present and calibrated with no quality issues; \'Suspect\': at least one spectrum is missing or calibrated with quality issues; \'Failed\': no calibrated spectra." ;
		:qa_pct_data_missing = 100.f ;
		:qa_pct_data_geo = 0.f ;
		:qa_pct_data_sci_mode = 0.f ;
		string :qa_no_data = "TRUE" ;
		string :title = "13:30 orbit L1 CHIRP" ;
		string :summary = "The CHIRP Level 1 product for the 13:30 sun-synchronous orbit consists of calibrated radiance spectra at a common resolution derived from hyperspectral instruments on EOS-Aqua, S-NPP, and JPSS-1/NOAA-20 platforms adjusted to form a continuous climate-quality record." ;
		string :shortname = "SSYN1330CHIRP1_placeholder" ;
		string :product_group = "l1_chirp" ;
		string :metadata_link = "http://disc.sci.gsfc.nasa.gov/" ;
		string :references = "" ;
		string :contributor_name = "UMBC Atmospheric Spectroscopy Laboratory: Larrabee Strow" ;
		string :contributor_role = "CrIS L1B Scientist" ;
		:wnum_delta_lw = 0.625f ;
		:wnum_delta_mw = 0.8333333f ;
		:wnum_delta_sw = 1.25f ;
}
